`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    11:06:26 11/13/2022 
// Design Name: 
// Module Name:    MReg 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module MReg(
    input [1:0] WDSelE,
    input RFenE,
    input FWSelE,
	 input [1:0] BEmodE,
	 input [2:0] BEXTOpE,
    input [31:0] ALUOutE,
    input [31:0] RD2SE,
	 input [31:0] HLE,
    input [4:0] A1E,
    input [4:0] A2E,
    input [2:0] TnewE,
    input [4:0] A3E,
    input [31:0] PC8E,
    input clk,
	 input reset,
	 input Req,
    output [1:0] WDSelM,
    output RFenM,
    output FWSelM,
	 output [1:0] BEmodM,
	 output [2:0] BEXTOpM,
    output [31:0] ALUOutM,
    output [31:0] RD2SM,
	 output [31:0] HLM,
    output [4:0] A1M,
    output [4:0] A2M,
    output [2:0] TnewM,
	 output [4:0] A3M,
    output [31:0] PC8M,
	 input [4:0] ExcE,
	 output [4:0] ExcEM,
	 input BDInE,
	 output BDInM,
	 input MTC0E,
	 output MTC0M,
	 input ERETE,
	 output ERETM,
	 input [4:0] ACP0E,
	 output [4:0] ACP0M
    );
	reg [1:0] WDSelreg;
   reg RFenreg;
   reg FWSelreg;
	reg [1:0] BEmodreg;
	reg [2:0] BEXTOpreg;
   reg [31:0] ALUOutreg;
	reg [31:0] RD2Sreg;
	reg [31:0] HLreg;
   reg [4:0] A1reg;
   reg [4:0] A2reg;
   reg [2:0] Tnewreg;
   reg [4:0] A3reg;
   reg [31:0] PC8reg;
	reg [4:0] Excreg;
	reg BDInreg;
	reg MTC0reg;
	reg ERETreg;
	reg [4:0] ACP0reg;
	initial begin
		WDSelreg <= 2'd0;
		RFenreg <= 1'd0;
		FWSelreg <= 1'd0;
		BEmodreg <= 2'd0;
		BEXTOpreg <= 3'd0;
		ALUOutreg <= 32'd0;
		RD2Sreg <= 32'd0;
		HLreg <= 32'd0;
		A1reg <= 5'd0;
		A2reg <= 5'd0;
		Tnewreg <= 3'd0;
		A3reg <= 5'd0;
		PC8reg <= 32'h3000 + 32'd8;
		Excreg <= 5'd0;
		BDInreg <= 1'd0;
		MTC0reg <= 1'd0;
		ERETreg <= 1'd0;
		ACP0reg <= 5'd0;
	end
	always@(posedge clk)begin
		if(reset || Req)begin
			WDSelreg <= 2'd0;
			RFenreg <= 1'd0;
			FWSelreg <= 1'd0;
			BEmodreg <= 2'd0;
			BEXTOpreg <= 3'd0;
			ALUOutreg <= 32'd0;
			RD2Sreg <= 32'd0;
			HLreg <= 32'd0;
			A1reg <= 5'd0;
			A2reg <= 5'd0;
			Tnewreg <= 3'd0;
			A3reg <= 5'd0;
			PC8reg <= ((Req)? (32'h4180 + 32'd8) : (32'h3000 + 32'd8));
			Excreg <= 5'd0;
			BDInreg <= 1'd0;
			MTC0reg <= 1'd0;
			ERETreg <= 1'd0;
			ACP0reg <= 5'd0;
		end else begin
			WDSelreg <= WDSelE;
			RFenreg <= RFenE;
			FWSelreg <= FWSelE;
			BEmodreg <= BEmodE;
			BEXTOpreg <= BEXTOpE;
			ALUOutreg <= ALUOutE;
			RD2Sreg <= RD2SE;
			HLreg <= HLE;
			A1reg <= A1E;
			A2reg <= A2E;
			Tnewreg <= TnewE;
			A3reg <= A3E;
			PC8reg <= PC8E;
			Excreg <= ExcE;
			BDInreg <= BDInE;
			MTC0reg <= MTC0E;
			ERETreg <= ERETE;
			ACP0reg <= ACP0E;
		end
	end
	assign WDSelM = WDSelreg;
   assign RFenM = RFenreg;
   assign FWSelM = FWSelreg;
	assign BEmodM = BEmodreg;
	assign BEXTOpM = BEXTOpreg;
   assign ALUOutM = ALUOutreg;
	assign RD2SM = RD2Sreg;
	assign HLM = HLreg;
   assign A1M = A1reg;
   assign A2M = A2reg;
   assign TnewM = (Tnewreg == 0) ? 3'd0 : (Tnewreg - 1);
   assign A3M = A3reg;
   assign PC8M = PC8reg;
	assign ExcEM = Excreg;
	assign BDInM = BDInreg;
	assign MTC0M = MTC0reg;
	assign ERETM = ERETreg;
	assign ACP0M = ACP0reg;
endmodule
